
package body mypackage is
  constant five :integer := four +1;
end package body mypackage;
