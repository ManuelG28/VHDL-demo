library ieee;
use ieee.std_logic_1164.all;
use work.mypackage.all;

entity mymodule is
	port( clk: in std_logic
	);
end mymodule;

architecture sim of mymodule is
begin
	process
	 constant t:integer := four;
	begin
	
	end process;
end architecture sim;