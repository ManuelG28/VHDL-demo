
architecture rtl of mymodule is
begin
	process
	begin
	
	end process;
end architecture rtl;