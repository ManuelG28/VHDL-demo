
package mypackage is
   constant four :integer := 4;
end package mypackage;
